`timescale 1ns / 1ps

module singlecycle(
		   input	     reset, //Active High
		   input [63:0]	     startpc,
		   output reg [63:0] currentpc,
		   output [63:0]     MemtoRegOut, // this should be
						   // attached to the
						   // output of the
						   // MemtoReg Mux
		   input	     CLK
		   );

   // Next PC connections
   wire [63:0] 			     nextpc;       // The next PC, to be updated on clock cycle

   // Instruction Memory connections
   wire [31:0] 			     instruction;  // The current instruction

   // Parts of instruction
   wire [4:0] 			     rd;            // The destination register
   wire [4:0] 			     rm;            // Operand 1
   wire [4:0] 			     rn;            // Operand 2
   wire [10:0] 			     opcode;

   // Control wires
   wire 			     Reg2Loc;
   wire 			     ALUSrc;
   wire 			     MemtoReg;
   wire 			     RegWrite;
   wire 			     MemRead;
   wire 			     MemWrite;
   wire 			     Branch;
   wire 			     Uncondbranch;
   wire [3:0] 			     ALUop;
   wire [1:0] 			     SignOp;

   // Register file connections
   wire [63:0] 			     regoutA;     // Output A
   wire [63:0] 			     regoutB;     // Output B

   // ALU connections
   wire [63:0] 			     aluout;
   wire 			     zero;

   // Sign Extender connections
   wire [63:0] 			     extimm;

   // Data Memory connections
   wire [63:0]                       memout;

   // Multiplexer outputs
   wire [63:0]                       aluin2;      // ALU input 2 (from ALUSrc mux)

   // PC update logic
   always @(posedge CLK)
     begin
        if (reset)
          currentpc <= #3 startpc;
        else
          currentpc <= #3 nextpc;
     end

   // Debug output - use negedge to avoid race conditions
   always @(negedge CLK)
     begin
        if (currentpc >= 64'h0 && currentpc <= 64'h30)
          $display("  [negedge] PC=%h X9=%h X10=%h X11=%h X12=%h X13=%h BusA=%h BusB=%h ALUOut=%h",
                   currentpc, rf.rf[9], rf.rf[10], rf.rf[11], rf.rf[12], rf.rf[13], regoutA, regoutB, aluout);
     end

   // Parts of instruction
   assign rd = instruction[4:0];
   assign rm = instruction[9:5];
   assign rn = Reg2Loc ? instruction[4:0] : instruction[20:16];
   assign opcode = instruction[31:21];

   // Instruction Memory
   InstructionMemory imem(
			  .Data(instruction),
			  .Address(currentpc)
			  );





// get the instruction at current pc, then decompose into rd, rm, rn, opcode. [6] (in schematic)
// contorl unit input = opcode, output [2] (in schematic)






   // Control Unit
   SC_Control SingleCycleControl(
		   .Reg2Loc(Reg2Loc),
		   .ALUSrc(ALUSrc),
		   .MemtoReg(MemtoReg),
		   .RegWrite(RegWrite),
		   .MemRead(MemRead),
		   .MemWrite(MemWrite),
		   .Branch(Branch),
		   .Uncondbranch(Uncondbranch),
		   .ALUOp(ALUop),
		   .SignOp(SignOp),
		   .opcode(opcode)
		   );







// registerfile [2] and [5]
// output is BusA[read data 1] and BusB[read data2]



   // Register File
   RegisterFile rf(
		   .BusA(regoutA),
		   .BusB(regoutB),
		   .BusW(MemtoRegOut),
		   .RA(rm),
		   .RB(rn),
		   .RW(rd),
		   .RegWr(RegWrite),
		   .Clk(CLK)
		   );





// sign extend immediates so its 64 bits so u can add with other 64 bits such as registers 

   // Sign Extender
   SignExtender signext(
			.SignExOut(extimm),
			.Instruction(instruction),
			.SignOp(SignOp)
			);







// [2]
   // ALUSrc Multiplexer: selects between regoutB and sign-extended immediate
   assign aluin2 = ALUSrc ? extimm : regoutB;




// [6]
// input either BusA [read data 1] or BusB aluin2[2, a mux to select between extended immedaite or regout B]
   // ALU
   ALU alu(
	   .BusW(aluout),
	   .BusA(regoutA),
	   .BusB(aluin2),
	   .ALUCtrl(ALUop),
	   .Zero(zero)
	   );





//  memwrite and memread [blue] 
   // Data Memory
   DataMemory datamem(
		      .ReadData(memout),
		      .Address(aluout),
		      .WriteData(regoutB),
		      .MemoryRead(MemRead),
		      .MemoryWrite(MemWrite),
		      .Clock(CLK)
		      );

   // MemtoReg Multiplexer: selects between ALU output and memory output
   assign MemtoRegOut = MemtoReg ? memout : aluout;

   // Next PC Logic
   NextPClogic nextpclogic(
			   .NextPC(nextpc),
			   .CurrentPC(currentpc),
			   .SignExtImm64(extimm),
			   .Branch(Branch),
			   .ALUZero(zero),
			   .Uncondbranch(Uncondbranch)
			   );

endmodule
